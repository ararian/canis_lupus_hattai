

// デコーダ
module decoder(input logic pc, output xx);



endmodule


