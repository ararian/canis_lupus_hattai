
// //TODO:下記の命令を実装予定
// LB = 10'h003, 
// LH = 10'h083,
// LW = 10'h103, 
// LBU = 10'h203,
// LHU = 10'h283, 
