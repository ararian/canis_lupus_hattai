
// module writeback()

// ({decodeToExecOrDmem.next_funct3, decodeToExecOrDmem.next_opcode}) 

// endmodule