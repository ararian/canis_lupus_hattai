package defs;
    parameter MEM_SIZE = 4000-1;
endpackage
