
module writeback(
    execToWriteback.writeback execToWriteback, 
    dmemToWriteback.writeback dmemToWriteback
)

// ({decodeToExecOrDmem.next_funct3, decodeToExecOrDmem.next_opcode}) 

endmodule

